module ClockDivider (
    input wire clk,          // ����ʱ���ź�
    output wire sec_pulse    // ����������ź�
);

reg [24:0] counter = 0;     // �ڲ��Ĵ��������ڼ���ʱ������

always @(posedge clk) begin
    if (counter == 25000000) // ����ʹ��50 MHzʱ�ӣ�������25000000��ʾ1������
        counter <= 0;       // �����ﵽ���ֵ��λΪ0
    else
        counter <= counter + 1; // ��ÿ��ʱ���������Ӽ���ֵ
end

assign sec_pulse = (counter == 25000000); // �������ﵽ25000000ʱ������1������

endmodule
/*

�����ǽ���������ʱ���źŷ�ƵΪ1�������źš�
��ͨ��һ���ڲ��Ĵ��� counter ������ʱ�����ڣ��������ﵽ�ض�ֵ������50 MHzʱ����Ϊ25000000��ʱ��
����һ��1�������ź� sec_pulse�����ģ���������ͬ��������������ĳЩӦ������Ҫÿ�봥��һ�β���ʱ�ǳ����á�
*/