module CoinDetector (
    input wire [3:0] coin_input, // ����Ӳ���źţ����ڼ��Ӳ������
    output wire [3:0] coin_code  // ���Ӳ�ұ��룬��ʾ��⵽��Ӳ������
);

assign coin_code = coin_input; // ֱ�ӽ�Ӳ�������źŸ��Ƶ�Ӳ�ұ�������ź�

endmodule
/*

�����Ӳ���ź�ֱ�Ӹ��Ƶ�Ӳ�ұ�������źţ����ڽ�Ӳ��������Ϣ���ݸ�����ģ�顣
�����û�н����κ�Ӳ�����͵ļ������ת����ֻ�Ǽ򵥵ؽ������źŴ��ݵ�����˿ڣ�
�Թ�����ģ��ʹ�á����ģ����Ը��ݾ����Ӳ�Ҽ�����������չ��
*/